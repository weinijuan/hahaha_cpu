// `include "cpu.svh"
// module preif
//     import cpuDefine::*;
// #(
//     parameter WIDTH = 100
// ) (
//     input logic aclk,
//     input logic aresetn,
//     input logic valid_in,
//     input logic[WIDTH-1:0] data_in,
//     input logic ready_go,
//     input logic[WIDTH-1:0] nop_data,
//     input logic allow_in,
//     input logic flush,
//     output logic valid_out,
//     output logic[WIDTH-1:0] data_out,
//     output logic allow_out
// );

//     logic ready_go;
//     always_comb begin
//         if (ready_go) begin
//             data_out 
//         end
//     end
    



// endmodule
